module riscv(input clk, input reset)